module top(
    input ref_clk,
    output tmds_0_p,
    output tmds_0_n,
    output tmds_1_p,
    output tmds_1_n,
    output tmds_2_p,
    output tmds_2_n,
    output tmds_clk_p,
    output tmds_clk_n,
    output led_0,
    output led_1,
    output led_2,
    output led_3,
    output led_4
);


wire pxlclk_raw, pxlclk;
wire serclk_raw, serclk;
wire serclk_locked;
wire rstn;
reg [7:0] r, g, b;


SB_PLL40_CORE pll_serclk (
    .REFERENCECLK (ref_clk),
    .PLLOUTGLOBAL (serclk_raw),
    .LOCK (serclk_locked),
    .BYPASS (1'b0),
    .RESETB (1'b1)
);

defparam pll_serclk.FEEDBACK_PATH = "SIMPLE";
defparam pll_serclk.DIVR          = 4'b0000;
defparam pll_serclk.DIVF          = 7'b1010011;
defparam pll_serclk.DIVQ          = 3'b011;
defparam pll_serclk.FILTER_RANGE  = 3'b001;


SB_GB serclk_gb (
    .USER_SIGNAL_TO_GLOBAL_BUFFER (serclk_raw),
    .GLOBAL_BUFFER_OUTPUT (serclk)
);

clk_divider pxlclk_divider (
    .clki (serclk),
    .clko (pxlclk_raw)
);

SB_GB pxlclk_gb (
    .USER_SIGNAL_TO_GLOBAL_BUFFER (pxlclk_raw),
    .GLOBAL_BUFFER_OUTPUT (pxlclk)
);

assign rstn = serclk_locked;

reg [9:0] col_cnt;
reg [9:0] row_cnt;

reg hsync, vsync, dena;

initial begin
    r <= 8'b00000000;
    g <= 8'b00000000;
    b <= 8'b00000000;

    col_cnt <= 0;
    row_cnt <= 0;

    hsync <= 0;
    vsync <= 0;
    dena  <= 0;
end

always @(posedge pxlclk) begin
    
    col_cnt <= col_cnt + 1;
    if (col_cnt == 16-1) begin
    // hsync pulse
    hsync <= 1'b1;
    end else if (col_cnt == 112-1) begin
        // back porch
        hsync <= 1'b0;
    end else if (col_cnt == 160-1) begin
        dena <= 1'b1;
    end else if (col_cnt == 800-1) begin
        dena <= 1'b0;
        col_cnt <= 0;
        row_cnt <= row_cnt + 1;
    end

    if (row_cnt > 480-1) begin
        dena <= 1'b0;
        if (row_cnt == 490-1) begin
            vsync <= 1'b1;
        end else if (row_cnt == 492-1) begin
            vsync <= 1'b0;
        end else if (row_cnt == 525-1) begin
            row_cnt <= 0;
        end
    end

end


dvi tmds (
    .serclk (serclk),
    .pxlclk (pxlclk),
    .rstn   (rstn),
    .r      (r),
    .g      (g),
    .b      (b),
    .hsync  (hsync),
    .vsync  (vsync),
    .dena   (dena),
    .tmds_p ({tmds_clk_p, tmds_2_p, tmds_1_p, tmds_0_p}),
    .tmds_n ({tmds_clk_n, tmds_2_n, tmds_1_n, tmds_0_n})
);

assign led_0 = 0;
assign led_1 = 0;
assign led_2 = 0;
assign led_3 = 0;
assign led_4 = rstn;



wire [7:0] char_line;

character_generator cg_0 (
    .pxlclk (pxlclk),
	.ascii  (col_cnt[9:3]),
	.row    (row_cnt[2:0]),
	.dout   (char_line)
);

reg [2:0] char_col;
reg pxl;
always @(posedge pxlclk) begin
	pxl <= char_line[char_col];
	char_col <= char_col + 1;
	if (pxl) begin
		r <= 8'hFF;
		g <= 8'hFF;
		b <= 8'hFF;
	end else begin
		r <= 8'h00;
		g <= 8'h00;
		b <= 8'h00;
	end
end




endmodule
